module main

import mana

fn main() {
	mana.start()
}
