module main

import mana

fn main() {
	mana.start(2)
}
