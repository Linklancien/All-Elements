module main

import gg
import mana

const bg_color = gg.Color{0, 0, 0, 255}

struct App {
mut:
	ctx &gg.Context = unsafe { nil }

	player_pool mana.Mana_pool
}

fn main() {
	mut app := &App{}
	app.ctx = gg.new_context(
		width:        100 * 8
		height:       100 * 6
		window_title: '-Render Life-'
		user_data:    app
		bg_color:     bg_color
		frame_fn:     on_frame
		sample_count: 4
	)

	app.player_pool = mana.Mana_pool{
		elements_list:     [mana.Elements.water, mana.Elements.air, mana.Elements.fire,
			mana.Elements.earth]
		elements_quantity: [f32(1), 15, 25, 2]
	}

	app.ctx.run()
}

fn on_frame(mut app App) {
	app.ctx.begin()
	app.player_pool.render(400, 300, 50, 20, app.ctx)
	app.ctx.end()
}
